module den
  (
    input clk,
    input d,
    output dout
  );
  reg[16] data='b45;
  always @ (posedge clk)
  begin

    c/c++
    python
    c#
    





  end
endmodule
